module q7_14 (in, out);
    input [4;0] in;
    output [4:0] out;
endmodule